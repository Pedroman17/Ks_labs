library verilog;
use verilog.vl_types.all;
entity f4_1 is
    port(
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        f_1             : out    vl_logic
    );
end f4_1;
